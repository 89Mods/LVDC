module ttl_74ahc1g04(
	input a,
	output y
);

assign #4 y = !a;

endmodule
