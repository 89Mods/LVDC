module ttl_74hct32(
	input a1,
	input b1,
	output y1,
	input a2,
	input b2,
	output y2,
	input a3,
	input b3,
	output y3,
	input a4,
	input b4,
	output y4
);

assign #16 y1 = a1 | b1;
assign #16 y2 = a2 | b2;
assign #16 y3 = a3 | b3;
assign #16 y4 = a4 | b4;

endmodule
