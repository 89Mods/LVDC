module ttl_74lv1t34(
	input A,
	output Y
);

assign Y = A;

endmodule
